../mult16x9/deploy/csa.sv