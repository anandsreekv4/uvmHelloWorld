// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : afifo_tb
//
// File Name: afifo_read_sequencer.sv
//
//
// Version:   1.0
//
//=============================================================================
// Description: Sequencer for afifo_read
//=============================================================================

`ifndef AFIFO_READ_SEQUENCER_SV
`define AFIFO_READ_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(rd_transaction) afifo_read_sequencer_t;


`endif // AFIFO_READ_SEQUENCER_SV

