// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Copyright (c) Anand Sreekumar
//=============================================================================
// Project  : ../../design/afifo
//
// File Name: afifo_write_driver.sv
//
// Author   : Name   : Anand Sreekumar
//            Email  : anandsreekv4@gmail.com
//            Year   : 2021
//
// Version:   1.0
//
//=============================================================================
// Description: Driver for afifo_write
//=============================================================================

`ifndef AFIFO_WRITE_DRIVER_SV
`define AFIFO_WRITE_DRIVER_SV

// You can insert code here by setting driver_inc_before_class in file afifo_wr_if.tpl

class afifo_write_driver extends uvm_driver #(wr_transaction);

  `uvm_component_utils(afifo_write_driver)

  virtual afifo_write_if vif;

  afifo_write_config     m_config;

  extern function new(string name, uvm_component parent);

  // Methods run_phase and do_drive generated by setting driver_inc in file afifo_wr_if.tpl
  extern task run_phase(uvm_phase phase);
  extern task do_drive();

  // You can insert code here by setting driver_inc_inside_class in file afifo_wr_if.tpl

endclass : afifo_write_driver 


function afifo_write_driver::new(string name, uvm_component parent);
  super.new(name, parent);
endfunction : new


task afifo_write_driver::run_phase(uvm_phase phase);
  `uvm_info(get_type_name(), "run_phase", UVM_HIGH)

  forever
  begin
    seq_item_port.get_next_item(req);
      `uvm_info(get_type_name(), {"req item\n",req.sprint}, UVM_HIGH)
    do_drive();
    seq_item_port.item_done();
  end
endtask : run_phase


// Start of inlined include file ../../design/afifo/tb/include/afifo_write_do_drive.sv
task afifo_write_driver::do_drive();
    @(posedge vif.wclk_i);
    vif.winc_i <= req.winc; // modification so winc only when out of reset
    vif.wdata_i<= req.wdata;
    vif.wrstn_i<= req.wrstn;
    @(posedge vif.wclk_i);
    vif.winc_i <= 0;
endtask: do_drive
// End of inlined include file

// You can insert code here by setting driver_inc_after_class in file afifo_wr_if.tpl

`endif // AFIFO_WRITE_DRIVER_SV

