// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Copyright (c) Anand Sreekumar
//=============================================================================
// Project  : ../../design/afifo
//
// File Name: afifo_write_monitor.sv
//
// Author   : Name   : Anand Sreekumar
//            Email  : anandsreekv4@gmail.com
//            Year   : 2021
//
// Version:   1.0
//
//=============================================================================
// Description: Monitor for afifo_write
//=============================================================================

`ifndef AFIFO_WRITE_MONITOR_SV
`define AFIFO_WRITE_MONITOR_SV

// You can insert code here by setting monitor_inc_before_class in file afifo_wr_if.tpl

class afifo_write_monitor extends uvm_monitor;

  `uvm_component_utils(afifo_write_monitor)

  virtual afifo_write_if vif;

  afifo_write_config     m_config;

  uvm_analysis_port #(wr_transaction) analysis_port;

  wr_transaction m_trans;

  extern function new(string name, uvm_component parent);

  // Methods run_phase, and do_mon generated by setting monitor_inc in file afifo_wr_if.tpl
  extern task run_phase(uvm_phase phase);
  extern task do_mon();

  // You can insert code here by setting monitor_inc_inside_class in file afifo_wr_if.tpl

endclass : afifo_write_monitor 


function afifo_write_monitor::new(string name, uvm_component parent);
  super.new(name, parent);
  analysis_port = new("analysis_port", this);
endfunction : new


task afifo_write_monitor::run_phase(uvm_phase phase);
  `uvm_info(get_type_name(), "run_phase", UVM_HIGH)

  m_trans = wr_transaction::type_id::create("m_trans");
  do_mon();
endtask : run_phase


// Start of inlined include file ../../design/afifo/tb/include/afifo_write_do_mon.sv
task afifo_write_monitor::do_mon();
    string s;
    forever begin
        @(posedge vif.wclk_i);
        m_trans = wr_transaction::type_id::create("m_trans");
        m_trans.wdata = vif.wdata_i;
        m_trans.wrstn = vif.wrstn_i;
        m_trans.fifo_full = vif.fifo_full_o;
        m_trans.fifo_overflow = vif.fifo_ovflw_o;

        s = $sformatf("Sending following trn for coverage:-\n%s", m_trans.convert2string());
        `uvm_info(get_type_name(), s, UVM_DEBUG)
        analysis_port.write(m_trans);
    end
endtask: do_mon
// End of inlined include file

// You can insert code here by setting monitor_inc_after_class in file afifo_wr_if.tpl

`endif // AFIFO_WRITE_MONITOR_SV

