    // uvm_objection obj = phase.get_objection();
    // obj.set_drain_time(this, 1000ns);
    phase.phase_done.set_drain_time(this, 1000ns);
