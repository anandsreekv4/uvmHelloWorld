../mult16x9/deploy/fulladder.sv