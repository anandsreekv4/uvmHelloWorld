../mult16x9/deploy/mult_xy.sv