../mult16x9/deploy/mult16x9behav.sv