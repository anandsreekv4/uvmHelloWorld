// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : afifo_tb
//
// File Name: top_config.sv
//
//
// Version:   1.0
//
//=============================================================================
// Description: Configuration for top
//=============================================================================

`ifndef TOP_CONFIG_SV
`define TOP_CONFIG_SV

// You can insert code here by setting top_env_config_inc_before_class in file common.tpl

class top_config extends uvm_object;

  // Do not register config class with the factory

  virtual afifo_write_if   afifo_write_vif;            
  virtual afifo_read_if    afifo_read_vif;             

  uvm_active_passive_enum  is_active_afifo_write       = UVM_ACTIVE;
  uvm_active_passive_enum  is_active_afifo_read        = UVM_ACTIVE;

  bit                      checks_enable_afifo_write;  
  bit                      checks_enable_afifo_read;   

  bit                      coverage_enable_afifo_write;
  bit                      coverage_enable_afifo_read; 

  // You can insert variables here by setting config_var in file common.tpl

  // You can remove new by setting top_env_config_generate_methods_inside_class = no in file common.tpl

  extern function new(string name = "");

  // You can insert code here by setting top_env_config_inc_inside_class in file common.tpl

endclass : top_config 


// You can remove new by setting top_env_config_generate_methods_after_class = no in file common.tpl

function top_config::new(string name = "");
  super.new(name);

  // You can insert code here by setting top_env_config_append_to_new in file common.tpl

endfunction : new


// You can insert code here by setting top_env_config_inc_after_class in file common.tpl

`endif // TOP_CONFIG_SV

