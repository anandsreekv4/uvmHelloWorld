// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : afifo_tb
//
// File Name: afifo_read_monitor.sv
//
//
// Version:   1.0
//
//=============================================================================
// Description: Monitor for afifo_read
//=============================================================================

`ifndef AFIFO_READ_MONITOR_SV
`define AFIFO_READ_MONITOR_SV

// You can insert code here by setting monitor_inc_before_class in file afifo_rd_if.tpl

class afifo_read_monitor extends uvm_monitor;

  `uvm_component_utils(afifo_read_monitor)

  virtual afifo_read_if vif;

  afifo_read_config     m_config;

  uvm_analysis_port #(rd_transaction) analysis_port;

  rd_transaction m_trans;

  extern function new(string name, uvm_component parent);

  // Methods run_phase, and do_mon generated by setting monitor_inc in file afifo_rd_if.tpl
  extern task run_phase(uvm_phase phase);
  extern task do_mon();

  // You can insert code here by setting monitor_inc_inside_class in file afifo_rd_if.tpl

endclass : afifo_read_monitor 


function afifo_read_monitor::new(string name, uvm_component parent);
  super.new(name, parent);
  analysis_port = new("analysis_port", this);
endfunction : new


task afifo_read_monitor::run_phase(uvm_phase phase);
  `uvm_info(get_type_name(), "run_phase", UVM_HIGH)

  m_trans = rd_transaction::type_id::create("m_trans");
  do_mon();
endtask : run_phase


// Start of inlined include file afifo_tb/tb/include/afifo_read_do_mon.sv
task afifo_read_monitor::do_mon();
    string s;
    forever begin
        @(posedge vif.rclk_i);
        m_trans = rd_transaction::type_id::create("m_trans");
        m_trans.rdata = vif.rdata_o;
        m_trans.rrstn = vif.rrstn_i;
        m_trans.fifo_empty = vif.fifo_empty_o;
        m_trans.fifo_underflow = vif.fifo_undrflw_o;

        s = $sformatf("Sending following trn for coverage:-\n%s", m_trans.convert2string());
        `uvm_info(get_type_name(), s, UVM_MEDIUM)
        analysis_port.write(m_trans);
    end
endtask: do_mon
// End of inlined include file

// You can insert code here by setting monitor_inc_after_class in file afifo_rd_if.tpl

`endif // AFIFO_READ_MONITOR_SV

