../mult16x9/deploy/ppg.sv