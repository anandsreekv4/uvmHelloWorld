../mult16x9/deploy/cpa.sv